CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
149
13 Logic Switch~
5 370 1549 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3343 0 0
2
45171.8 0
0
13 Logic Switch~
5 250 1546 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7923 0 0
2
45171.8 0
0
13 Logic Switch~
5 273 1545 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6174 0 0
2
45171.8 44
0
13 Logic Switch~
5 298 1545 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6692 0 0
2
45171.8 43
0
13 Logic Switch~
5 320 1546 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8790 0 0
2
45171.8 42
0
13 Logic Switch~
5 394 1548 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4595 0 0
2
45171.8 41
0
13 Logic Switch~
5 415 1549 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
667 0 0
2
45171.8 40
0
13 Logic Switch~
5 435 1549 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8743 0 0
2
45171.8 39
0
13 Logic Switch~
5 382 532 0 10 11
0 91 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8298 0 0
2
45171.5 0
0
13 Logic Switch~
5 362 532 0 10 11
0 104 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
313 0 0
2
45171.5 0
0
13 Logic Switch~
5 341 531 0 10 11
0 120 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7548 0 0
2
45171.5 0
0
13 Logic Switch~
5 293 529 0 10 11
0 92 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8973 0 0
2
45171.5 0
0
13 Logic Switch~
5 270 529 0 10 11
0 103 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9712 0 0
2
45171.5 0
0
13 Logic Switch~
5 247 529 0 10 11
0 119 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4518 0 0
2
45171.5 0
0
13 Logic Switch~
5 252 161 0 10 11
0 122 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5596 0 0
2
5.90089e-315 0
0
13 Logic Switch~
5 251 297 0 10 11
0 123 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
692 0 0
2
5.90089e-315 0
0
13 Logic Switch~
5 251 256 0 10 11
0 124 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6258 0 0
2
5.90089e-315 0
0
13 Logic Switch~
5 251 210 0 10 11
0 121 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5578 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 867 2983 0 3 22
0 14 13 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 37 0
1 U
8709 0 0
2
45171.9 5
0
9 2-In AND~
219 868 3033 0 3 22
0 13 12 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 34 0
1 U
9131 0 0
2
45171.9 4
0
9 2-In AND~
219 866 2935 0 3 22
0 14 12 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 34 0
1 U
3645 0 0
2
45171.9 3
0
6 74136~
219 857 2869 0 3 22
0 13 14 26
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU6B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 36 0
1 U
7613 0 0
2
45171.9 2
0
6 74136~
219 935 2902 0 3 22
0 26 12 11
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU6A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 36 0
1 U
9467 0 0
2
45171.9 1
0
8 3-In OR~
219 971 2988 0 4 22
0 25 24 23 10
0
0 0 624 0
4 4075
-14 -24 14 -16
6 CARR1A
-13 -25 29 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 35 0
1 U
3932 0 0
2
45171.9 0
0
9 2-In AND~
219 974 2719 0 3 22
0 18 22 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 34 0
1 U
5288 0 0
2
45171.9 5
0
9 2-In AND~
219 975 2769 0 3 22
0 17 22 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
4934 0 0
2
45171.9 4
0
9 2-In AND~
219 973 2671 0 3 22
0 18 17 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
5987 0 0
2
45171.9 3
0
6 74136~
219 964 2605 0 3 22
0 17 22 30
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU5D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 33 0
1 U
7737 0 0
2
45171.9 2
0
6 74136~
219 1042 2638 0 3 22
0 30 18 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 33 0
1 U
4200 0 0
2
45171.9 1
0
8 3-In OR~
219 1078 2724 0 4 22
0 29 28 27 12
0
0 0 624 0
4 4075
-14 -24 14 -16
6 CARR3C
-13 -25 29 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 31 0
1 U
5780 0 0
2
45171.9 0
0
8 3-In OR~
219 803 2727 0 4 22
0 33 32 31 13
0
0 0 624 0
4 4075
-14 -24 14 -16
6 CARR3A
-13 -25 29 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 31 0
1 U
6490 0 0
2
45171.9 5
0
6 74136~
219 767 2641 0 3 22
0 34 20 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUD
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
8663 0 0
2
45171.9 4
0
6 74136~
219 689 2608 0 3 22
0 19 21 34
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUC
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
318 0 0
2
45171.9 3
0
9 2-In AND~
219 698 2674 0 3 22
0 20 19 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 29 0
1 U
348 0 0
2
45171.9 2
0
9 2-In AND~
219 700 2772 0 3 22
0 21 19 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
8551 0 0
2
45171.9 1
0
9 2-In AND~
219 699 2722 0 3 22
0 21 20 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 29 0
1 U
7295 0 0
2
45171.9 0
0
8 3-In OR~
219 1226 2467 0 4 22
0 40 39 38 18
0
0 0 624 0
4 4075
-14 -24 14 -16
5 CARRY
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 24 0
1 U
9900 0 0
2
45171.9 5
0
6 74136~
219 1190 2381 0 3 22
0 41 37 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
8725 0 0
2
45171.9 4
0
6 74136~
219 1112 2348 0 3 22
0 35 36 41
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU4A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
366 0 0
2
45171.9 3
0
9 2-In AND~
219 1121 2414 0 3 22
0 37 36 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
5762 0 0
2
45171.9 2
0
9 2-In AND~
219 1123 2512 0 3 22
0 36 35 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
4943 0 0
2
45171.9 1
0
9 2-In AND~
219 1122 2462 0 3 22
0 37 35 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
3435 0 0
2
45171.9 0
0
8 3-In OR~
219 966 2468 0 4 22
0 47 46 45 20
0
0 0 624 0
4 4075
-14 -24 14 -16
6 CARR2B
-13 -25 29 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 24 0
1 U
8705 0 0
2
45171.9 5
0
6 74136~
219 930 2382 0 3 22
0 48 43 36
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U10C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
4331 0 0
2
45171.9 4
0
6 74136~
219 852 2349 0 3 22
0 42 44 48
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U10D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
787 0 0
2
45171.9 3
0
9 2-In AND~
219 861 2415 0 3 22
0 44 42 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
3655 0 0
2
45171.9 2
0
9 2-In AND~
219 863 2513 0 3 22
0 42 43 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
6682 0 0
2
45171.9 1
0
9 2-In AND~
219 862 2463 0 3 22
0 44 43 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
582 0 0
2
45171.9 0
0
6 74136~
219 668 2378 0 3 22
0 49 50 44
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U10B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 27 0
1 U
3125 0 0
2
45171.9 0
0
9 2-In AND~
219 542 2476 0 3 22
0 4 5 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A2B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
5466 0 0
2
45171.9 0
0
9 2-In AND~
219 542 2545 0 3 22
0 6 3 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B3
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
52 0 0
2
45171.9 0
0
9 2-In AND~
219 543 2886 0 3 22
0 2 3 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A3B3
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
3898 0 0
2
45171.9 0
0
9 2-In AND~
219 545 2628 0 3 22
0 2 5 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A3B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 25 0
1 U
9413 0 0
2
45171.9 0
0
9 2-In AND~
219 545 2802 0 3 22
0 4 3 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A2B3
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 25 0
1 U
8576 0 0
2
45171.9 0
0
9 2-In AND~
219 677 2435 0 3 22
0 50 49 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
622 0 0
2
45171.9 0
0
9 2-In AND~
219 542 2375 0 3 22
0 2 7 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A3B1
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
9152 0 0
2
45171.9 0
0
6 74136~
219 1165 2078 0 3 22
0 51 52 53
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 22 0
1 U
783 0 0
2
45171.9 0
0
9 2-In AND~
219 1175 2146 0 3 22
0 51 52 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 23 0
1 U
4262 0 0
2
45171.9 0
0
8 3-In OR~
219 1022 2157 0 4 22
0 59 58 57 43
0
0 0 624 0
4 4075
-14 -24 14 -16
6 CARR2A
-13 -25 29 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 24 0
1 U
6121 0 0
2
45171.9 5
0
9 2-In AND~
219 942 2167 0 3 22
0 54 56 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
3879 0 0
2
45171.9 4
0
9 2-In AND~
219 943 2216 0 3 22
0 55 56 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0BD
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
7345 0 0
2
45171.9 3
0
9 2-In AND~
219 942 2120 0 3 22
0 55 54 59
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0BC
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
3198 0 0
2
45171.9 2
0
6 74136~
219 1024 2073 0 3 22
0 56 60 51
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU3B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
9849 0 0
2
45171.9 1
0
6 74136~
219 936 2060 0 3 22
0 55 54 60
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU3A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
479 0 0
2
45171.9 0
0
8 3-In OR~
219 761 2140 0 4 22
0 66 65 64 49
0
0 0 624 0
4 4075
-14 -24 14 -16
5 carry
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 12 0
1 U
3905 0 0
2
45171.9 5
0
9 2-In AND~
219 681 2150 0 3 22
0 63 61 65
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
4394 0 0
2
45171.9 4
0
9 2-In AND~
219 682 2199 0 3 22
0 62 61 64
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
4391 0 0
2
45171.9 3
0
9 2-In AND~
219 681 2103 0 3 22
0 63 62 66
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
3681 0 0
2
45171.9 2
0
6 74136~
219 763 2056 0 3 22
0 63 67 55
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 sum
-7 -27 14 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
6466 0 0
2
45171.9 1
0
6 74136~
219 673 2045 0 3 22
0 62 61 67
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU1C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
5230 0 0
2
45171.9 0
0
9 2-In AND~
219 545 2229 0 3 22
0 6 5 54
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 23 0
1 U
8324 0 0
2
45171.9 0
0
14 Logic Display~
6 1102 1543 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3445 0 0
2
45171.8 0
0
14 Logic Display~
6 1151 1545 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7543 0 0
2
45171.8 0
0
9 2-In AND~
219 536 1602 0 3 22
0 8 9 81
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B0
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
6187 0 0
2
45171.8 38
0
9 2-In AND~
219 537 1664 0 3 22
0 6 9 80
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B0
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
5476 0 0
2
45171.8 37
0
9 2-In AND~
219 537 1790 0 3 22
0 9 4 75
0
0 0 624 0
0
4 A2B0
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
3936 0 0
2
45171.8 36
0
9 2-In AND~
219 538 1710 0 3 22
0 8 7 79
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
5770 0 0
2
45171.8 35
0
9 2-In AND~
219 540 1869 0 3 22
0 6 7 76
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
7884 0 0
2
45171.8 34
0
9 2-In AND~
219 545 1957 0 3 22
0 8 5 70
0
0 0 624 0
4 A0B2
-14 -24 14 -16
4 A0B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
3690 0 0
2
45171.8 33
0
9 2-In AND~
219 546 2051 0 3 22
0 2 9 61
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A3B0
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
3611 0 0
2
45171.8 32
0
9 2-In AND~
219 547 2120 0 3 22
0 4 7 62
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A2B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
7912 0 0
2
45171.8 31
0
9 2-In AND~
219 544 2282 0 3 22
0 8 3 52
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B3
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
6416 0 0
2
45171.8 30
0
14 Logic Display~
6 1229 1545 0 1 2
10 68
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7278 0 0
2
45171.8 29
0
14 Logic Display~
6 1177 1545 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6804 0 0
2
45171.8 28
0
14 Logic Display~
6 1201 1545 0 1 2
10 53
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9568 0 0
2
45171.8 27
0
14 Logic Display~
6 1279 1545 0 1 2
10 81
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7178 0 0
2
45171.8 26
0
14 Logic Display~
6 1254 1543 0 1 2
10 78
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7982 0 0
2
45171.8 25
0
14 Logic Display~
6 1128 1545 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
513 0 0
2
45171.8 24
0
6 74136~
219 681 1646 0 3 22
0 79 80 78
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
8190 0 0
2
45171.8 23
0
9 2-In AND~
219 688 1696 0 3 22
0 80 79 74
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-18 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
5209 0 0
2
45171.8 22
0
6 74136~
219 677 1771 0 3 22
0 76 75 77
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 SU2C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
7239 0 0
2
45171.8 21
0
6 74136~
219 782 1774 0 3 22
0 74 77 69
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 sum
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
9474 0 0
2
45171.8 20
0
9 2-In AND~
219 684 1816 0 3 22
0 75 76 73
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
3783 0 0
2
45171.8 19
0
9 2-In AND~
219 685 1860 0 3 22
0 74 76 72
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
5422 0 0
2
45171.8 18
0
9 2-In AND~
219 687 1907 0 3 22
0 75 74 71
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
8527 0 0
2
45171.8 17
0
8 3-In OR~
219 779 1838 0 4 22
0 73 71 72 63
0
0 0 624 0
4 4075
-14 -24 14 -16
5 carry
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 12 0
1 U
761 0 0
2
45171.8 16
0
6 74136~
219 929 1779 0 3 22
0 69 70 68
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
7323 0 0
2
45171.8 15
0
9 2-In AND~
219 937 1837 0 3 22
0 70 69 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
8543 0 0
2
45171.8 14
0
8 3-In OR~
219 719 1312 0 4 22
0 86 85 84 82
0
0 0 624 0
4 4075
-14 -24 14 -16
5 CARRY
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 8 0
1 U
4240 0 0
2
45171.8 0
0
6 74136~
219 683 1226 0 3 22
0 87 88 83
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7857 0 0
2
45171.8 0
0
6 74136~
219 605 1193 0 3 22
0 89 90 87
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUB
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7255 0 0
2
45171.8 0
0
8 3-In OR~
219 868 1109 0 4 22
0 95 94 93 88
0
0 0 624 0
4 4075
-14 -24 14 -16
5 CARRY
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 8 0
1 U
7736 0 0
2
45171.8 0
0
9 2-In AND~
219 614 1259 0 3 22
0 90 89 86
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
5435 0 0
2
45171.8 0
0
9 2-In AND~
219 616 1357 0 3 22
0 89 88 84
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3446 0 0
2
45171.8 0
0
9 2-In AND~
219 788 1119 0 3 22
0 98 96 94
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3914 0 0
2
45171.8 0
0
9 2-In AND~
219 789 1168 0 3 22
0 97 96 93
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3948 0 0
2
45171.8 0
0
9 2-In AND~
219 615 1307 0 3 22
0 90 88 85
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3901 0 0
2
45171.8 0
0
9 2-In AND~
219 788 1072 0 3 22
0 97 98 95
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
6295 0 0
2
45171.8 0
0
9 2-In AND~
219 622 1094 0 3 22
0 102 101 89
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 carry
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
332 0 0
2
45171.8 0
0
6 74136~
219 870 1025 0 3 22
0 96 99 100
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9737 0 0
2
45171.8 0
0
6 74136~
219 780 1014 0 3 22
0 97 98 99
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUD
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
9910 0 0
2
45171.8 0
0
6 74136~
219 618 1032 0 3 22
0 102 101 98
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 sum
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3834 0 0
2
45171.8 0
0
9 2-In AND~
219 884 820 0 3 22
0 107 106 96
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3138 0 0
2
45171.8 0
0
6 74136~
219 876 762 0 3 22
0 106 107 105
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
5409 0 0
2
45171.8 0
0
8 3-In OR~
219 726 821 0 4 22
0 110 108 109 102
0
0 0 624 0
4 4075
-14 -24 14 -16
5 carry
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
983 0 0
2
45171.8 0
0
9 2-In AND~
219 634 890 0 3 22
0 112 111 108
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6652 0 0
2
45171.8 0
0
9 2-In AND~
219 632 843 0 3 22
0 111 113 109
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4281 0 0
2
45171.8 0
0
9 2-In AND~
219 631 799 0 3 22
0 112 113 110
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
6847 0 0
2
45171.8 0
0
6 74136~
219 729 757 0 3 22
0 111 114 106
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 sum
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6543 0 0
2
45171.8 0
0
6 74136~
219 624 754 0 3 22
0 113 112 114
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUD
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7168 0 0
2
45171.8 0
0
9 2-In AND~
219 635 679 0 3 22
0 117 116 111
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-18 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3828 0 0
2
45171.8 0
0
6 74136~
219 628 629 0 3 22
0 116 117 115
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
955 0 0
2
45171.8 0
0
14 Logic Display~
6 863 537 0 1 2
10 82
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7782 0 0
2
45171.6 0
0
14 Logic Display~
6 980 536 0 1 2
10 115
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
824 0 0
2
45171.6 0
0
14 Logic Display~
6 1009 534 0 1 2
10 118
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6983 0 0
2
45171.6 0
0
14 Logic Display~
6 921 537 0 1 2
10 100
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3185 0 0
2
45171.6 0
0
14 Logic Display~
6 893 537 0 1 2
10 83
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4213 0 0
2
45171.6 0
0
14 Logic Display~
6 949 537 0 1 2
10 105
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 P2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9765 0 0
2
45171.6 0
0
9 2-In AND~
219 490 1237 0 3 22
0 92 91 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A2B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8986 0 0
2
45171.6 0
0
9 2-In AND~
219 494 1103 0 3 22
0 91 103 97
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3273 0 0
2
45171.6 0
0
9 2-In AND~
219 493 1034 0 3 22
0 92 104 101
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A2B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5636 0 0
2
45171.6 0
0
9 2-In AND~
219 492 940 0 3 22
0 119 91 107
0
0 0 624 0
4 A0B2
-14 -24 14 -16
4 A0B2
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
327 0 0
2
45171.6 0
0
9 2-In AND~
219 487 852 0 3 22
0 104 103 113
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9233 0 0
2
45171.6 0
0
9 2-In AND~
219 485 693 0 3 22
0 119 104 116
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3875 0 0
2
45171.6 0
0
9 2-In AND~
219 487 783 0 3 22
0 92 120 112
0
0 0 624 0
0
4 A2B0
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9991 0 0
2
45171.6 0
0
9 2-In AND~
219 484 647 0 3 22
0 103 120 117
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B0
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3221 0 0
2
45171.6 0
0
9 2-In AND~
219 483 585 0 3 22
0 120 119 118
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B0
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8874 0 0
2
45171.6 0
0
14 Logic Display~
6 738 347 0 1 2
10 125
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7400 0 0
2
5.90089e-315 0
0
14 Logic Display~
6 739 284 0 1 2
10 126
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3623 0 0
2
5.90089e-315 0
0
14 Logic Display~
6 738 224 0 1 2
10 127
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3311 0 0
2
5.90089e-315 0
0
14 Logic Display~
6 737 167 0 1 2
10 128
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5736 0 0
2
5.90089e-315 0
0
6 74136~
219 616 319 0 3 22
0 129 130 126
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3143 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 624 370 0 3 22
0 130 129 125
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5835 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 528 301 0 3 22
0 132 131 129
0
0 0 624 0
6 74LS08
-21 -24 21 -16
5 CARRY
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5108 0 0
2
5.90089e-315 0
0
6 74136~
219 520 251 0 3 22
0 131 132 127
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUM
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3320 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 401 348 0 3 22
0 123 121 130
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
523 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 401 293 0 3 22
0 122 123 132
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B1
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3557 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 401 235 0 3 22
0 121 124 131
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A1B0
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7246 0 0
2
5.90089e-315 0
0
9 2-In AND~
219 401 179 0 3 22
0 122 124 128
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 A0B0
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3916 0 0
2
5.90089e-315 0
0
258
0 1 2 0 0 8192 0 0 52 7 0 4
513 2619
506 2619
506 2877
519 2877
0 2 3 0 0 4096 0 0 52 3 0 3
501 2811
501 2895
519 2895
0 2 3 0 0 4096 0 0 54 8 0 3
481 2554
481 2811
521 2811
0 1 4 0 0 4096 0 0 54 11 0 3
491 2467
491 2793
521 2793
0 0 5 0 0 4096 0 0 0 15 6 2
504 2238
503 2485
2 2 5 0 0 16 0 53 50 0 0 4
521 2637
500 2637
500 2485
518 2485
1 1 2 0 0 0 0 56 53 0 0 4
518 2366
513 2366
513 2619
521 2619
0 2 3 0 0 4096 0 0 51 10 0 3
457 2291
457 2554
518 2554
0 1 6 0 0 4096 0 0 51 16 0 3
467 2220
467 2536
518 2536
1 2 3 0 0 4224 0 8 82 0 0 3
435 1561
435 2291
520 2291
0 1 4 0 0 4224 0 0 50 18 0 3
476 2111
476 2467
518 2467
0 2 7 0 0 4096 0 0 56 17 0 3
497 2129
497 2384
518 2384
0 1 2 0 0 4096 0 0 56 21 0 3
488 2042
488 2366
518 2366
0 1 8 0 0 4224 0 0 82 139 0 3
353 1593
353 2273
520 2273
0 2 5 0 0 4096 0 0 71 128 0 3
504 1966
504 2238
521 2238
0 1 6 0 0 4224 0 0 71 137 0 3
380 1655
380 2220
521 2220
0 2 7 0 0 4224 0 0 81 134 0 3
429 1719
429 2129
523 2129
0 1 4 0 0 0 0 0 81 133 0 3
448 1799
448 2111
523 2111
2 0 9 0 0 4096 0 80 0 0 20 2
522 2060
464 2060
0 2 9 0 0 4224 0 0 80 138 0 3
464 1611
464 2060
522 2060
1 1 2 0 0 4224 0 5 80 0 0 3
320 1558
320 2042
522 2042
0 4 10 0 0 16384 0 0 24 23 0 6
1401 2342
1404 2342
1404 2364
1405 2364
1405 2988
1004 2988
1 0 10 0 0 12416 0 72 0 0 22 5
1102 1561
1102 1623
1401 1623
1401 2346
1404 2346
1 3 11 0 0 12416 0 88 23 0 0 7
1128 1563
1128 1612
1380 1612
1380 2329
1378 2329
1378 2902
968 2902
0 2 12 0 0 8192 0 0 20 26 0 4
811 2944
813 2944
813 3042
844 3042
0 2 12 0 0 0 0 0 21 32 0 6
900 2885
894 2885
894 2901
811 2901
811 2944
842 2944
2 0 13 0 0 4096 0 19 0 0 28 4
843 2992
831 2992
831 2993
826 2993
0 1 13 0 0 8320 0 0 20 33 0 4
840 2830
826 2830
826 3024
844 3024
0 1 14 0 0 8192 0 0 19 30 0 4
831 2924
835 2924
835 2974
843 2974
0 1 14 0 0 0 0 0 21 31 0 3
831 2886
831 2926
842 2926
3 2 14 0 0 4224 0 52 22 0 0 4
564 2886
833 2886
833 2878
841 2878
4 2 12 0 0 12416 0 30 23 0 0 6
1111 2724
1115 2724
1115 2814
900 2814
900 2911
919 2911
4 1 13 0 0 0 0 31 22 0 0 6
836 2727
840 2727
840 2850
836 2850
836 2860
841 2860
1 3 15 0 0 20608 0 73 29 0 0 7
1151 1563
1151 1585
1311 1585
1311 2059
1312 2059
1312 2638
1075 2638
1 3 16 0 0 12416 0 84 38 0 0 5
1177 1563
1177 1573
1297 1573
1297 2381
1223 2381
0 1 17 0 0 4096 0 0 26 37 0 3
881 2680
881 2760
951 2760
2 0 17 0 0 0 0 27 0 0 41 3
949 2680
879 2680
879 2641
0 1 18 0 0 8192 0 0 25 39 0 4
926 2660
927 2660
927 2710
950 2710
0 1 18 0 0 4096 0 0 27 40 0 4
1006 2647
926 2647
926 2662
949 2662
4 2 18 0 0 12416 0 37 29 0 0 6
1259 2467
1263 2467
1263 2555
1006 2555
1006 2647
1026 2647
3 1 17 0 0 4224 0 32 28 0 0 4
800 2641
935 2641
935 2596
948 2596
0 2 19 0 0 8192 0 0 35 43 0 4
642 2683
644 2683
644 2781
676 2781
0 2 19 0 0 0 0 0 34 49 0 4
665 2595
642 2595
642 2683
674 2683
0 2 20 0 0 4096 0 0 36 45 0 3
656 2665
656 2731
675 2731
0 1 20 0 0 4096 0 0 34 48 0 4
736 2641
656 2641
656 2665
674 2665
0 1 21 0 0 8192 0 0 35 47 0 4
664 2713
668 2713
668 2763
676 2763
0 1 21 0 0 4096 0 0 36 50 0 3
664 2628
664 2713
675 2713
4 2 20 0 0 12416 0 43 32 0 0 8
999 2468
1003 2468
1003 2537
736 2537
736 2661
743 2661
743 2650
751 2650
3 1 19 0 0 16512 0 55 33 0 0 6
698 2435
726 2435
726 2463
665 2463
665 2599
673 2599
3 2 21 0 0 4224 0 53 33 0 0 4
566 2628
665 2628
665 2617
673 2617
2 0 22 0 0 8192 0 25 0 0 53 3
950 2728
950 2730
940 2730
2 0 22 0 0 4096 0 26 0 0 53 2
951 2778
940 2778
3 2 22 0 0 4224 0 54 28 0 0 4
566 2802
940 2802
940 2614
948 2614
3 3 23 0 0 4224 0 20 24 0 0 4
889 3033
950 3033
950 2997
958 2997
3 2 24 0 0 4224 0 19 24 0 0 4
888 2983
950 2983
950 2988
959 2988
3 1 25 0 0 4224 0 21 24 0 0 4
887 2935
950 2935
950 2979
958 2979
3 1 26 0 0 8320 0 22 23 0 0 4
890 2869
911 2869
911 2893
919 2893
3 3 27 0 0 4224 0 26 30 0 0 4
996 2769
1057 2769
1057 2733
1065 2733
3 2 28 0 0 4224 0 25 30 0 0 4
995 2719
1057 2719
1057 2724
1066 2724
3 1 29 0 0 4224 0 27 30 0 0 4
994 2671
1057 2671
1057 2715
1065 2715
3 1 30 0 0 8320 0 28 29 0 0 4
997 2605
1018 2605
1018 2629
1026 2629
3 3 31 0 0 4224 0 35 31 0 0 4
721 2772
782 2772
782 2736
790 2736
3 2 32 0 0 4224 0 36 31 0 0 4
720 2722
782 2722
782 2727
791 2727
3 1 33 0 0 4224 0 34 31 0 0 4
719 2674
782 2674
782 2718
790 2718
3 1 34 0 0 8320 0 33 32 0 0 4
722 2608
743 2608
743 2632
751 2632
1 0 35 0 0 8192 0 39 0 0 68 3
1096 2339
1026 2339
1026 2545
2 2 35 0 0 0 0 42 41 0 0 4
1098 2471
1086 2471
1086 2521
1099 2521
3 2 35 0 0 4224 0 51 41 0 0 4
563 2545
1091 2545
1091 2521
1099 2521
0 1 36 0 0 8320 0 0 41 70 0 4
1073 2423
1091 2423
1091 2503
1099 2503
0 2 36 0 0 0 0 0 40 78 0 3
1073 2392
1073 2423
1097 2423
0 1 37 0 0 8192 0 0 42 72 0 4
1089 2404
1085 2404
1085 2453
1098 2453
0 1 37 0 0 4096 0 0 40 73 0 4
1159 2380
1089 2380
1089 2405
1097 2405
3 2 37 0 0 16512 0 58 38 0 0 6
1196 2146
1235 2146
1235 2181
1159 2181
1159 2390
1174 2390
3 3 38 0 0 4224 0 41 37 0 0 4
1144 2512
1205 2512
1205 2476
1213 2476
3 2 39 0 0 4224 0 42 37 0 0 4
1143 2462
1205 2462
1205 2467
1214 2467
3 1 40 0 0 4224 0 40 37 0 0 4
1142 2414
1205 2414
1205 2458
1213 2458
3 1 41 0 0 8320 0 39 38 0 0 4
1145 2348
1166 2348
1166 2372
1174 2372
3 2 36 0 0 0 0 44 39 0 0 6
963 2382
1018 2382
1018 2392
1083 2392
1083 2357
1096 2357
1 0 42 0 0 8192 0 45 0 0 80 4
836 2340
817 2340
817 2424
818 2424
0 2 42 0 0 0 0 0 46 81 0 3
818 2476
818 2424
837 2424
3 1 42 0 0 4224 0 50 47 0 0 4
563 2476
823 2476
823 2504
839 2504
4 2 43 0 0 12416 0 59 44 0 0 6
1055 2157
1059 2157
1059 2247
901 2247
901 2391
914 2391
3 0 44 0 0 4096 0 49 0 0 92 3
701 2378
761 2378
761 2393
3 3 45 0 0 4224 0 47 43 0 0 4
884 2513
945 2513
945 2477
953 2477
3 2 46 0 0 4224 0 48 43 0 0 4
883 2463
945 2463
945 2468
954 2468
3 1 47 0 0 4224 0 46 43 0 0 4
882 2415
945 2415
945 2459
953 2459
3 1 48 0 0 8320 0 45 44 0 0 4
885 2349
906 2349
906 2373
914 2373
0 2 43 0 0 0 0 0 47 89 0 3
831 2483
831 2522
839 2522
0 2 43 0 0 0 0 0 48 82 0 7
907 2391
907 2402
908 2402
908 2483
830 2483
830 2472
838 2472
0 1 44 0 0 0 0 0 48 91 0 4
828 2406
825 2406
825 2454
838 2454
0 1 44 0 0 0 0 0 46 92 0 3
828 2393
828 2406
837 2406
3 2 44 0 0 4224 0 0 45 0 0 4
758 2393
828 2393
828 2358
836 2358
0 2 49 0 0 4096 0 0 55 95 0 3
648 2369
648 2444
653 2444
0 1 50 0 0 8192 0 0 55 96 0 4
637 2385
638 2385
638 2426
653 2426
4 1 49 0 0 12416 0 65 49 0 0 6
794 2140
798 2140
798 2224
644 2224
644 2369
652 2369
3 2 50 0 0 4224 0 56 49 0 0 4
563 2375
637 2375
637 2387
652 2387
0 1 51 0 0 4096 0 0 58 98 0 3
1116 2073
1116 2137
1151 2137
3 1 51 0 0 4224 0 63 57 0 0 4
1057 2073
1141 2073
1141 2069
1149 2069
2 0 52 0 0 8192 0 57 0 0 100 4
1149 2087
1140 2087
1140 2159
1143 2159
3 2 52 0 0 4224 0 82 58 0 0 4
565 2282
1143 2282
1143 2155
1151 2155
1 3 53 0 0 4224 0 85 57 0 0 3
1201 1563
1201 2078
1198 2078
3 0 54 0 0 4224 0 71 0 0 114 4
566 2229
899 2229
899 2080
904 2080
0 1 55 0 0 8192 0 0 61 104 0 4
877 2108
878 2108
878 2207
919 2207
0 1 55 0 0 0 0 0 62 105 0 3
877 2056
877 2111
918 2111
3 1 55 0 0 4224 0 69 64 0 0 4
796 2056
907 2056
907 2051
920 2051
3 0 56 0 0 8192 0 98 0 0 111 3
958 1837
962 1837
962 2027
3 3 57 0 0 8320 0 61 59 0 0 4
964 2216
996 2216
996 2166
1009 2166
3 2 58 0 0 12416 0 60 59 0 0 4
963 2167
983 2167
983 2157
1010 2157
3 1 59 0 0 4224 0 62 59 0 0 4
963 2120
1001 2120
1001 2148
1009 2148
2 0 56 0 0 0 0 60 0 0 111 2
918 2176
914 2176
2 1 56 0 0 8320 0 61 63 0 0 8
919 2225
914 2225
914 2027
1002 2027
1002 2039
1000 2039
1000 2064
1008 2064
0 1 54 0 0 0 0 0 60 114 0 3
907 2129
907 2158
918 2158
3 2 60 0 0 4224 0 64 63 0 0 4
969 2060
992 2060
992 2082
1008 2082
2 2 54 0 0 0 0 62 64 0 0 6
918 2129
904 2129
904 2080
910 2080
910 2069
920 2069
0 2 61 0 0 4096 0 0 67 116 0 3
635 2159
635 2208
658 2208
0 2 61 0 0 4224 0 0 66 123 0 3
615 2051
615 2159
657 2159
0 1 62 0 0 8192 0 0 67 118 0 4
636 2120
645 2120
645 2190
658 2190
0 2 62 0 0 0 0 0 68 122 0 3
636 2120
636 2112
657 2112
0 1 63 0 0 8192 0 0 66 120 0 4
644 2094
649 2094
649 2141
657 2141
0 1 63 0 0 8192 0 0 68 121 0 4
739 1975
644 1975
644 2094
657 2094
4 1 63 0 0 16512 0 96 69 0 0 6
812 1838
816 1838
816 1920
739 1920
739 2047
747 2047
3 1 62 0 0 8320 0 81 70 0 0 4
568 2120
639 2120
639 2036
657 2036
3 2 61 0 0 0 0 80 70 0 0 4
567 2051
649 2051
649 2054
657 2054
3 3 64 0 0 8320 0 67 65 0 0 4
703 2199
735 2199
735 2149
748 2149
3 2 65 0 0 12416 0 66 65 0 0 4
702 2150
722 2150
722 2140
749 2140
3 1 66 0 0 4224 0 68 65 0 0 4
702 2103
740 2103
740 2131
748 2131
3 2 67 0 0 4224 0 70 69 0 0 4
706 2045
731 2045
731 2065
747 2065
1 2 5 0 0 4224 0 7 79 0 0 3
415 1561
415 1966
521 1966
1 1 8 0 0 0 0 77 79 0 0 4
514 1701
498 1701
498 1948
521 1948
0 2 7 0 0 0 0 0 78 134 0 3
494 1719
494 1878
516 1878
0 1 6 0 0 0 0 0 78 137 0 3
481 1655
481 1860
516 1860
0 1 9 0 0 0 0 0 76 136 0 5
506 1673
506 1770
505 1770
505 1781
513 1781
2 1 4 0 0 0 0 76 4 0 0 3
513 1799
298 1799
298 1557
1 2 7 0 0 0 0 6 77 0 0 3
394 1560
394 1719
514 1719
0 1 8 0 0 0 0 0 77 139 0 3
493 1593
493 1701
514 1701
0 2 9 0 0 0 0 0 75 138 0 3
506 1611
506 1673
513 1673
1 1 6 0 0 0 0 3 75 0 0 3
273 1557
273 1655
513 1655
1 2 9 0 0 0 0 1 74 0 0 3
370 1561
370 1611
512 1611
1 1 8 0 0 0 0 2 74 0 0 3
250 1558
250 1593
512 1593
3 1 68 0 0 4224 0 97 83 0 0 3
962 1779
1229 1779
1229 1563
0 2 69 0 0 4224 0 0 98 144 0 3
876 1762
876 1846
913 1846
1 0 70 0 0 4096 0 98 0 0 143 2
913 1828
905 1828
3 2 70 0 0 4224 0 79 97 0 0 4
566 1957
905 1957
905 1788
913 1788
3 1 69 0 0 0 0 92 97 0 0 6
815 1774
876 1774
876 1762
905 1762
905 1770
913 1770
3 2 71 0 0 8320 0 95 96 0 0 4
708 1907
753 1907
753 1838
767 1838
3 3 72 0 0 4224 0 94 96 0 0 4
706 1860
758 1860
758 1847
766 1847
3 1 73 0 0 4224 0 93 96 0 0 4
705 1816
758 1816
758 1829
766 1829
1 2 74 0 0 8192 0 94 95 0 0 4
661 1851
645 1851
645 1916
663 1916
0 2 74 0 0 4224 0 0 95 156 0 5
722 1696
722 1927
655 1927
655 1916
663 1916
0 1 75 0 0 4224 0 0 95 155 0 3
640 1800
640 1898
663 1898
0 2 76 0 0 4096 0 0 94 154 0 2
648 1869
661 1869
1 0 75 0 0 0 0 93 0 0 155 3
660 1807
660 1800
653 1800
2 0 76 0 0 0 0 93 0 0 154 2
660 1825
648 1825
3 1 76 0 0 8320 0 78 91 0 0 4
561 1869
648 1869
648 1762
661 1762
3 2 75 0 0 0 0 76 91 0 0 6
558 1790
640 1790
640 1800
653 1800
653 1780
661 1780
3 1 74 0 0 0 0 90 92 0 0 4
709 1696
726 1696
726 1765
766 1765
3 2 77 0 0 12416 0 91 92 0 0 4
710 1771
725 1771
725 1783
766 1783
3 1 78 0 0 4224 0 89 87 0 0 3
714 1646
1254 1646
1254 1561
1 0 79 0 0 8192 0 89 0 0 160 3
665 1637
634 1637
634 1710
3 2 79 0 0 4224 0 77 90 0 0 4
559 1710
656 1710
656 1705
664 1705
0 1 80 0 0 4096 0 0 90 162 0 3
656 1664
656 1687
664 1687
3 2 80 0 0 4224 0 75 89 0 0 4
558 1664
657 1664
657 1655
665 1655
3 1 81 0 0 4224 0 74 86 0 0 3
557 1602
1279 1602
1279 1563
4 1 82 0 0 8320 0 99 123 0 0 5
752 1312
967 1312
967 575
863 575
863 555
3 1 83 0 0 8320 0 100 127 0 0 5
716 1226
938 1226
938 563
893 563
893 555
3 3 84 0 0 4224 0 104 99 0 0 4
637 1357
698 1357
698 1321
706 1321
3 2 85 0 0 4224 0 107 99 0 0 4
636 1307
698 1307
698 1312
707 1312
3 1 86 0 0 4224 0 103 99 0 0 4
635 1259
698 1259
698 1303
706 1303
3 1 87 0 0 8320 0 101 100 0 0 4
638 1193
659 1193
659 1217
667 1217
0 2 88 0 0 4096 0 0 104 171 0 3
579 1327
579 1366
592 1366
0 2 88 0 0 8192 0 0 107 172 0 5
661 1246
661 1327
578 1327
578 1316
591 1316
4 2 88 0 0 12416 0 102 100 0 0 6
901 1109
905 1109
905 1246
659 1246
659 1235
667 1235
0 1 89 0 0 8192 0 0 104 174 0 4
572 1268
584 1268
584 1348
592 1348
0 2 89 0 0 8320 0 0 103 178 0 4
581 1171
572 1171
572 1268
590 1268
0 1 90 0 0 8192 0 0 107 176 0 4
581 1250
578 1250
578 1298
591 1298
0 1 90 0 0 0 0 0 103 177 0 3
581 1237
581 1250
590 1250
3 2 90 0 0 4224 0 129 101 0 0 4
511 1237
581 1237
581 1202
589 1202
3 1 89 0 0 0 0 109 101 0 0 6
643 1094
647 1094
647 1161
581 1161
581 1184
589 1184
0 2 91 0 0 4096 0 0 129 200 0 3
463 1094
463 1246
466 1246
0 1 92 0 0 8192 0 0 129 202 0 4
428 1022
453 1022
453 1228
466 1228
3 3 93 0 0 8320 0 106 102 0 0 4
810 1168
842 1168
842 1118
855 1118
3 2 94 0 0 12416 0 105 102 0 0 4
809 1119
829 1119
829 1109
856 1109
3 1 95 0 0 4224 0 108 102 0 0 4
809 1072
847 1072
847 1100
855 1100
2 0 96 0 0 4096 0 105 0 0 185 2
764 1128
760 1128
2 0 96 0 0 8320 0 106 0 0 191 5
765 1177
760 1177
760 979
848 979
848 991
0 1 97 0 0 4096 0 0 106 189 0 3
737 1063
737 1159
765 1159
0 1 98 0 0 4096 0 0 105 188 0 3
753 1081
753 1110
764 1110
0 2 98 0 0 4096 0 0 108 193 0 3
750 1032
750 1081
764 1081
0 1 97 0 0 0 0 0 108 192 0 3
737 1000
737 1063
764 1063
3 2 99 0 0 4224 0 111 110 0 0 4
813 1014
838 1014
838 1034
854 1034
3 1 96 0 0 0 0 113 110 0 0 6
905 820
909 820
909 991
848 991
848 1016
854 1016
3 1 97 0 0 12416 0 130 111 0 0 5
515 1103
558 1103
558 1000
764 1000
764 1005
3 2 98 0 0 4224 0 112 111 0 0 4
651 1032
756 1032
756 1023
764 1023
1 3 100 0 0 4224 0 126 110 0 0 3
921 555
921 1025
903 1025
0 2 101 0 0 4096 0 0 109 196 0 3
575 1034
575 1103
598 1103
3 2 101 0 0 4224 0 131 112 0 0 4
514 1034
594 1034
594 1041
602 1041
0 1 102 0 0 8192 0 0 109 198 0 4
594 1023
590 1023
590 1085
598 1085
4 1 102 0 0 12416 0 115 112 0 0 6
759 821
758 821
758 920
594 920
594 1023
602 1023
0 2 103 0 0 4224 0 0 130 229 0 3
437 861
437 1112
470 1112
0 1 91 0 0 0 0 0 130 227 0 3
446 949
446 1094
470 1094
0 2 104 0 0 4224 0 0 131 230 0 3
458 843
458 1043
469 1043
0 1 92 0 0 4224 0 0 131 232 0 3
428 774
428 1025
469 1025
3 1 105 0 0 8320 0 114 128 0 0 3
909 762
949 762
949 555
0 2 106 0 0 4224 0 0 113 207 0 3
823 745
823 829
860 829
1 0 107 0 0 4096 0 113 0 0 206 2
860 811
852 811
3 2 107 0 0 4224 0 132 114 0 0 4
513 940
852 940
852 771
860 771
3 1 106 0 0 0 0 119 114 0 0 6
762 757
823 757
823 745
852 745
852 753
860 753
3 2 108 0 0 8320 0 116 115 0 0 4
655 890
700 890
700 821
714 821
3 3 109 0 0 4224 0 117 115 0 0 4
653 843
705 843
705 830
713 830
3 1 110 0 0 4224 0 118 115 0 0 4
652 799
705 799
705 812
713 812
1 2 111 0 0 8192 0 117 116 0 0 4
608 834
592 834
592 899
610 899
0 2 111 0 0 4224 0 0 116 219 0 5
669 679
669 910
602 910
602 899
610 899
0 1 112 0 0 4224 0 0 116 218 0 3
587 783
587 881
610 881
0 2 113 0 0 4096 0 0 117 217 0 2
595 852
608 852
1 0 112 0 0 0 0 118 0 0 218 3
607 790
607 783
600 783
2 0 113 0 0 0 0 118 0 0 217 2
607 808
595 808
3 1 113 0 0 8320 0 133 120 0 0 4
508 852
595 852
595 745
608 745
3 2 112 0 0 0 0 135 120 0 0 4
508 783
600 783
600 763
608 763
3 1 111 0 0 0 0 121 119 0 0 4
656 679
673 679
673 748
713 748
3 2 114 0 0 12416 0 120 119 0 0 4
657 754
672 754
672 766
713 766
3 1 115 0 0 4224 0 122 124 0 0 3
661 629
980 629
980 554
1 0 116 0 0 8192 0 122 0 0 223 3
612 620
581 620
581 693
3 2 116 0 0 4224 0 134 121 0 0 4
506 693
603 693
603 688
611 688
0 1 117 0 0 4096 0 0 121 225 0 3
603 647
603 670
611 670
3 2 117 0 0 4224 0 136 122 0 0 4
505 647
604 647
604 638
612 638
3 1 118 0 0 4224 0 137 125 0 0 3
504 585
1009 585
1009 552
1 2 91 0 0 4224 0 9 132 0 0 3
382 544
382 949
468 949
0 1 119 0 0 4224 0 0 132 234 0 3
447 684
447 931
468 931
0 2 103 0 0 0 0 0 133 236 0 3
404 638
404 861
463 861
0 1 104 0 0 0 0 0 133 233 0 3
436 702
436 843
463 843
0 2 120 0 0 8320 0 0 135 235 0 4
449 656
454 656
454 792
463 792
1 1 92 0 0 0 0 12 135 0 0 3
293 541
293 774
463 774
1 2 104 0 0 0 0 10 134 0 0 3
362 544
362 702
461 702
0 1 119 0 0 0 0 0 134 237 0 3
439 594
439 684
461 684
0 2 120 0 0 0 0 0 136 238 0 3
449 576
449 656
460 656
1 1 103 0 0 0 0 13 136 0 0 3
270 541
270 638
460 638
1 2 119 0 0 0 0 14 137 0 0 3
247 541
247 594
459 594
1 1 120 0 0 0 0 11 137 0 0 3
341 543
341 576
459 576
0 2 121 0 0 4224 0 0 146 245 0 3
338 210
338 357
377 357
0 1 122 0 0 4224 0 0 147 246 0 3
352 161
352 284
377 284
0 1 123 0 0 4096 0 0 146 242 0 3
369 302
369 339
377 339
1 2 123 0 0 4224 0 16 147 0 0 4
263 297
369 297
369 302
377 302
2 2 124 0 0 8192 0 148 149 0 0 4
377 244
364 244
364 188
377 188
1 2 124 0 0 4224 0 17 148 0 0 4
263 256
369 256
369 244
377 244
1 1 121 0 0 0 0 18 148 0 0 4
263 210
369 210
369 226
377 226
1 1 122 0 0 0 0 15 149 0 0 4
264 161
369 161
369 170
377 170
3 1 125 0 0 4224 0 143 138 0 0 3
645 370
738 370
738 365
3 1 126 0 0 4224 0 142 139 0 0 3
649 319
739 319
739 302
3 1 127 0 0 4224 0 145 140 0 0 3
553 251
738 251
738 242
3 1 128 0 0 4224 0 149 141 0 0 5
422 179
725 179
725 193
737 193
737 185
0 2 129 0 0 4224 0 0 143 254 0 3
577 301
577 379
600 379
2 1 130 0 0 8192 0 142 143 0 0 4
600 328
592 328
592 361
600 361
1 3 130 0 0 4224 0 143 146 0 0 4
600 361
430 361
430 348
422 348
3 1 129 0 0 0 0 144 142 0 0 4
549 301
592 301
592 310
600 310
0 2 131 0 0 4224 0 0 144 258 0 3
473 235
473 310
504 310
0 1 132 0 0 8192 0 0 144 257 0 3
495 293
495 292
504 292
3 2 132 0 0 4224 0 147 145 0 0 4
422 293
496 293
496 260
504 260
3 1 131 0 0 0 0 148 145 0 0 4
422 235
496 235
496 242
504 242
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
514 1479 661 1501
523 1486 651 1502
16 4 Bit Multiplier
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
461 462 600 486
466 466 594 482
16 3 Bit Multiplier
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
451 80 592 104
461 88 581 104
15 2 Bit Multipler
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
